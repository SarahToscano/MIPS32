module somasub_tb(a,b,cin,cout,s);

endmodule